-- Laboratory RA solutions/versuch4
-- Sommersemester 25
-- Group Details
-- Lab Date:
-- 1. Participant First and Last Name: 
-- 2. Participant First and Last Name:

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;
  use ieee.math_real.all;
  use work.constant_package.all;
  use work.types.all;

entity register_file is
-- begin solution:
   -- end solution!!
end entity register_file;

architecture behavior_debug of register_file is
-- begin solution:
   -- end solution!!
end architecture ;